VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_simple_riscv
  CLASS BLOCK ;
  FOREIGN tt_um_simple_riscv ;
  ORIGIN 0.000 0.000 ;
  SIZE 1440.320 BY 325.360 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 22.180 3.620 23.780 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 61.050 3.620 62.650 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 99.920 3.620 101.520 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 138.790 3.620 140.390 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 177.660 3.620 179.260 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 216.530 3.620 218.130 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 255.400 3.620 257.000 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 294.270 3.620 295.870 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 333.140 3.620 334.740 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 372.010 3.620 373.610 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 410.880 3.620 412.480 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 449.750 3.620 451.350 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 488.620 3.620 490.220 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 527.490 3.620 529.090 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 566.360 3.620 567.960 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 605.230 3.620 606.830 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 644.100 3.620 645.700 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 682.970 3.620 684.570 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 721.840 3.620 723.440 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 760.710 3.620 762.310 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 799.580 3.620 801.180 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 838.450 3.620 840.050 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 877.320 3.620 878.920 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 916.190 3.620 917.790 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 955.060 3.620 956.660 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 993.930 3.620 995.530 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1032.800 3.620 1034.400 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1071.670 3.620 1073.270 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1110.540 3.620 1112.140 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1149.410 3.620 1151.010 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1188.280 3.620 1189.880 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1227.150 3.620 1228.750 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1266.020 3.620 1267.620 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1304.890 3.620 1306.490 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1343.760 3.620 1345.360 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1382.630 3.620 1384.230 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1421.500 3.620 1423.100 321.740 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 18.880 3.620 20.480 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 57.750 3.620 59.350 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 96.620 3.620 98.220 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 135.490 3.620 137.090 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 174.360 3.620 175.960 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 213.230 3.620 214.830 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.100 3.620 253.700 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 290.970 3.620 292.570 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.840 3.620 331.440 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 368.710 3.620 370.310 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 407.580 3.620 409.180 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 446.450 3.620 448.050 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 485.320 3.620 486.920 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 524.190 3.620 525.790 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 563.060 3.620 564.660 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 601.930 3.620 603.530 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 640.800 3.620 642.400 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 679.670 3.620 681.270 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 718.540 3.620 720.140 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 757.410 3.620 759.010 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 796.280 3.620 797.880 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 835.150 3.620 836.750 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 874.020 3.620 875.620 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 912.890 3.620 914.490 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 951.760 3.620 953.360 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 990.630 3.620 992.230 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1029.500 3.620 1031.100 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1068.370 3.620 1069.970 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1107.240 3.620 1108.840 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1146.110 3.620 1147.710 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1184.980 3.620 1186.580 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1223.850 3.620 1225.450 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1262.720 3.620 1264.320 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1301.590 3.620 1303.190 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1340.460 3.620 1342.060 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1379.330 3.620 1380.930 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1418.200 3.620 1419.800 321.740 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    PORT
      LAYER Metal4 ;
        RECT 331.090 324.360 331.390 325.360 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 338.370 324.360 338.670 325.360 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    PORT
      LAYER Metal4 ;
        RECT 323.810 324.360 324.110 325.360 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    PORT
      LAYER Metal4 ;
        RECT 316.530 324.360 316.830 325.360 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    PORT
      LAYER Metal4 ;
        RECT 309.250 324.360 309.550 325.360 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    PORT
      LAYER Metal4 ;
        RECT 301.970 324.360 302.270 325.360 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    PORT
      LAYER Metal4 ;
        RECT 294.690 324.360 294.990 325.360 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    PORT
      LAYER Metal4 ;
        RECT 287.410 324.360 287.710 325.360 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    PORT
      LAYER Metal4 ;
        RECT 280.130 324.360 280.430 325.360 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    PORT
      LAYER Metal4 ;
        RECT 272.850 324.360 273.150 325.360 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    PORT
      LAYER Metal4 ;
        RECT 265.570 324.360 265.870 325.360 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    PORT
      LAYER Metal4 ;
        RECT 258.290 324.360 258.590 325.360 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 11.020000 ;
    PORT
      LAYER Metal4 ;
        RECT 251.010 324.360 251.310 325.360 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 243.730 324.360 244.030 325.360 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 236.450 324.360 236.750 325.360 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 229.170 324.360 229.470 325.360 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 221.890 324.360 222.190 325.360 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 214.610 324.360 214.910 325.360 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 207.330 324.360 207.630 325.360 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 83.570 324.360 83.870 325.360 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 76.290 324.360 76.590 325.360 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 69.010 324.360 69.310 325.360 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 61.730 324.360 62.030 325.360 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 54.450 324.360 54.750 325.360 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 47.170 324.360 47.470 325.360 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 39.890 324.360 40.190 325.360 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 32.610 324.360 32.910 325.360 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 141.810 324.360 142.110 325.360 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 134.530 324.360 134.830 325.360 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 127.250 324.360 127.550 325.360 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 119.970 324.360 120.270 325.360 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 112.690 324.360 112.990 325.360 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 105.410 324.360 105.710 325.360 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 98.130 324.360 98.430 325.360 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 90.850 324.360 91.150 325.360 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.604400 ;
    PORT
      LAYER Metal4 ;
        RECT 200.050 324.360 200.350 325.360 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.604400 ;
    PORT
      LAYER Metal4 ;
        RECT 192.770 324.360 193.070 325.360 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.604400 ;
    PORT
      LAYER Metal4 ;
        RECT 185.490 324.360 185.790 325.360 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.604400 ;
    PORT
      LAYER Metal4 ;
        RECT 178.210 324.360 178.510 325.360 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.604400 ;
    PORT
      LAYER Metal4 ;
        RECT 170.930 324.360 171.230 325.360 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.604400 ;
    PORT
      LAYER Metal4 ;
        RECT 163.650 324.360 163.950 325.360 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.604400 ;
    PORT
      LAYER Metal4 ;
        RECT 156.370 324.360 156.670 325.360 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.604400 ;
    PORT
      LAYER Metal4 ;
        RECT 149.090 324.360 149.390 325.360 ;
    END
  END uo_out[7]
  OBS
      LAYER Nwell ;
        RECT 2.930 319.280 1437.390 321.870 ;
      LAYER Pwell ;
        RECT 2.930 315.760 1437.390 319.280 ;
      LAYER Nwell ;
        RECT 2.930 311.440 1437.390 315.760 ;
      LAYER Pwell ;
        RECT 2.930 307.920 1437.390 311.440 ;
      LAYER Nwell ;
        RECT 2.930 303.600 1437.390 307.920 ;
      LAYER Pwell ;
        RECT 2.930 300.080 1437.390 303.600 ;
      LAYER Nwell ;
        RECT 2.930 295.760 1437.390 300.080 ;
      LAYER Pwell ;
        RECT 2.930 292.240 1437.390 295.760 ;
      LAYER Nwell ;
        RECT 2.930 287.920 1437.390 292.240 ;
      LAYER Pwell ;
        RECT 2.930 284.400 1437.390 287.920 ;
      LAYER Nwell ;
        RECT 2.930 280.080 1437.390 284.400 ;
      LAYER Pwell ;
        RECT 2.930 276.560 1437.390 280.080 ;
      LAYER Nwell ;
        RECT 2.930 272.240 1437.390 276.560 ;
      LAYER Pwell ;
        RECT 2.930 268.720 1437.390 272.240 ;
      LAYER Nwell ;
        RECT 2.930 264.400 1437.390 268.720 ;
      LAYER Pwell ;
        RECT 2.930 260.880 1437.390 264.400 ;
      LAYER Nwell ;
        RECT 2.930 256.560 1437.390 260.880 ;
      LAYER Pwell ;
        RECT 2.930 253.040 1437.390 256.560 ;
      LAYER Nwell ;
        RECT 2.930 248.720 1437.390 253.040 ;
      LAYER Pwell ;
        RECT 2.930 245.200 1437.390 248.720 ;
      LAYER Nwell ;
        RECT 2.930 240.880 1437.390 245.200 ;
      LAYER Pwell ;
        RECT 2.930 237.360 1437.390 240.880 ;
      LAYER Nwell ;
        RECT 2.930 233.040 1437.390 237.360 ;
      LAYER Pwell ;
        RECT 2.930 229.520 1437.390 233.040 ;
      LAYER Nwell ;
        RECT 2.930 225.200 1437.390 229.520 ;
      LAYER Pwell ;
        RECT 2.930 221.680 1437.390 225.200 ;
      LAYER Nwell ;
        RECT 2.930 217.360 1437.390 221.680 ;
      LAYER Pwell ;
        RECT 2.930 213.840 1437.390 217.360 ;
      LAYER Nwell ;
        RECT 2.930 209.520 1437.390 213.840 ;
      LAYER Pwell ;
        RECT 2.930 206.000 1437.390 209.520 ;
      LAYER Nwell ;
        RECT 2.930 201.680 1437.390 206.000 ;
      LAYER Pwell ;
        RECT 2.930 198.160 1437.390 201.680 ;
      LAYER Nwell ;
        RECT 2.930 193.840 1437.390 198.160 ;
      LAYER Pwell ;
        RECT 2.930 190.320 1437.390 193.840 ;
      LAYER Nwell ;
        RECT 2.930 186.000 1437.390 190.320 ;
      LAYER Pwell ;
        RECT 2.930 182.480 1437.390 186.000 ;
      LAYER Nwell ;
        RECT 2.930 178.160 1437.390 182.480 ;
      LAYER Pwell ;
        RECT 2.930 174.640 1437.390 178.160 ;
      LAYER Nwell ;
        RECT 2.930 170.320 1437.390 174.640 ;
      LAYER Pwell ;
        RECT 2.930 166.800 1437.390 170.320 ;
      LAYER Nwell ;
        RECT 2.930 162.480 1437.390 166.800 ;
      LAYER Pwell ;
        RECT 2.930 158.960 1437.390 162.480 ;
      LAYER Nwell ;
        RECT 2.930 154.640 1437.390 158.960 ;
      LAYER Pwell ;
        RECT 2.930 151.120 1437.390 154.640 ;
      LAYER Nwell ;
        RECT 2.930 146.800 1437.390 151.120 ;
      LAYER Pwell ;
        RECT 2.930 143.280 1437.390 146.800 ;
      LAYER Nwell ;
        RECT 2.930 138.960 1437.390 143.280 ;
      LAYER Pwell ;
        RECT 2.930 135.440 1437.390 138.960 ;
      LAYER Nwell ;
        RECT 2.930 131.120 1437.390 135.440 ;
      LAYER Pwell ;
        RECT 2.930 127.600 1437.390 131.120 ;
      LAYER Nwell ;
        RECT 2.930 123.280 1437.390 127.600 ;
      LAYER Pwell ;
        RECT 2.930 119.760 1437.390 123.280 ;
      LAYER Nwell ;
        RECT 2.930 115.440 1437.390 119.760 ;
      LAYER Pwell ;
        RECT 2.930 111.920 1437.390 115.440 ;
      LAYER Nwell ;
        RECT 2.930 107.600 1437.390 111.920 ;
      LAYER Pwell ;
        RECT 2.930 104.080 1437.390 107.600 ;
      LAYER Nwell ;
        RECT 2.930 99.760 1437.390 104.080 ;
      LAYER Pwell ;
        RECT 2.930 96.240 1437.390 99.760 ;
      LAYER Nwell ;
        RECT 2.930 91.920 1437.390 96.240 ;
      LAYER Pwell ;
        RECT 2.930 88.400 1437.390 91.920 ;
      LAYER Nwell ;
        RECT 2.930 84.080 1437.390 88.400 ;
      LAYER Pwell ;
        RECT 2.930 80.560 1437.390 84.080 ;
      LAYER Nwell ;
        RECT 2.930 76.240 1437.390 80.560 ;
      LAYER Pwell ;
        RECT 2.930 72.720 1437.390 76.240 ;
      LAYER Nwell ;
        RECT 2.930 68.400 1437.390 72.720 ;
      LAYER Pwell ;
        RECT 2.930 64.880 1437.390 68.400 ;
      LAYER Nwell ;
        RECT 2.930 60.560 1437.390 64.880 ;
      LAYER Pwell ;
        RECT 2.930 57.040 1437.390 60.560 ;
      LAYER Nwell ;
        RECT 2.930 52.720 1437.390 57.040 ;
      LAYER Pwell ;
        RECT 2.930 49.200 1437.390 52.720 ;
      LAYER Nwell ;
        RECT 2.930 44.880 1437.390 49.200 ;
      LAYER Pwell ;
        RECT 2.930 41.360 1437.390 44.880 ;
      LAYER Nwell ;
        RECT 2.930 37.040 1437.390 41.360 ;
      LAYER Pwell ;
        RECT 2.930 33.520 1437.390 37.040 ;
      LAYER Nwell ;
        RECT 2.930 29.200 1437.390 33.520 ;
      LAYER Pwell ;
        RECT 2.930 25.680 1437.390 29.200 ;
      LAYER Nwell ;
        RECT 2.930 21.360 1437.390 25.680 ;
      LAYER Pwell ;
        RECT 2.930 17.840 1437.390 21.360 ;
      LAYER Nwell ;
        RECT 2.930 13.520 1437.390 17.840 ;
      LAYER Pwell ;
        RECT 2.930 10.000 1437.390 13.520 ;
      LAYER Nwell ;
        RECT 2.930 5.680 1437.390 10.000 ;
      LAYER Pwell ;
        RECT 2.930 3.490 1437.390 5.680 ;
      LAYER Metal1 ;
        RECT 3.360 3.620 1436.960 321.740 ;
      LAYER Metal2 ;
        RECT 4.060 0.090 1422.960 325.270 ;
      LAYER Metal3 ;
        RECT 4.010 0.140 1423.010 325.220 ;
      LAYER Metal4 ;
        RECT 15.260 324.060 32.310 325.270 ;
        RECT 33.210 324.060 39.590 325.270 ;
        RECT 40.490 324.060 46.870 325.270 ;
        RECT 47.770 324.060 54.150 325.270 ;
        RECT 55.050 324.060 61.430 325.270 ;
        RECT 62.330 324.060 68.710 325.270 ;
        RECT 69.610 324.060 75.990 325.270 ;
        RECT 76.890 324.060 83.270 325.270 ;
        RECT 84.170 324.060 90.550 325.270 ;
        RECT 91.450 324.060 97.830 325.270 ;
        RECT 98.730 324.060 105.110 325.270 ;
        RECT 106.010 324.060 112.390 325.270 ;
        RECT 113.290 324.060 119.670 325.270 ;
        RECT 120.570 324.060 126.950 325.270 ;
        RECT 127.850 324.060 134.230 325.270 ;
        RECT 135.130 324.060 141.510 325.270 ;
        RECT 142.410 324.060 148.790 325.270 ;
        RECT 149.690 324.060 156.070 325.270 ;
        RECT 156.970 324.060 163.350 325.270 ;
        RECT 164.250 324.060 170.630 325.270 ;
        RECT 171.530 324.060 177.910 325.270 ;
        RECT 178.810 324.060 185.190 325.270 ;
        RECT 186.090 324.060 192.470 325.270 ;
        RECT 193.370 324.060 199.750 325.270 ;
        RECT 200.650 324.060 207.030 325.270 ;
        RECT 207.930 324.060 214.310 325.270 ;
        RECT 215.210 324.060 221.590 325.270 ;
        RECT 222.490 324.060 228.870 325.270 ;
        RECT 229.770 324.060 236.150 325.270 ;
        RECT 237.050 324.060 243.430 325.270 ;
        RECT 244.330 324.060 250.710 325.270 ;
        RECT 251.610 324.060 257.990 325.270 ;
        RECT 258.890 324.060 265.270 325.270 ;
        RECT 266.170 324.060 272.550 325.270 ;
        RECT 273.450 324.060 279.830 325.270 ;
        RECT 280.730 324.060 287.110 325.270 ;
        RECT 288.010 324.060 294.390 325.270 ;
        RECT 295.290 324.060 301.670 325.270 ;
        RECT 302.570 324.060 308.950 325.270 ;
        RECT 309.850 324.060 316.230 325.270 ;
        RECT 317.130 324.060 323.510 325.270 ;
        RECT 324.410 324.060 330.790 325.270 ;
        RECT 331.690 324.060 338.070 325.270 ;
        RECT 338.970 324.060 1371.300 325.270 ;
        RECT 15.260 322.040 1371.300 324.060 ;
        RECT 15.260 3.320 18.580 322.040 ;
        RECT 20.780 3.320 21.880 322.040 ;
        RECT 24.080 3.320 57.450 322.040 ;
        RECT 59.650 3.320 60.750 322.040 ;
        RECT 62.950 3.320 96.320 322.040 ;
        RECT 98.520 3.320 99.620 322.040 ;
        RECT 101.820 3.320 135.190 322.040 ;
        RECT 137.390 3.320 138.490 322.040 ;
        RECT 140.690 3.320 174.060 322.040 ;
        RECT 176.260 3.320 177.360 322.040 ;
        RECT 179.560 3.320 212.930 322.040 ;
        RECT 215.130 3.320 216.230 322.040 ;
        RECT 218.430 3.320 251.800 322.040 ;
        RECT 254.000 3.320 255.100 322.040 ;
        RECT 257.300 3.320 290.670 322.040 ;
        RECT 292.870 3.320 293.970 322.040 ;
        RECT 296.170 3.320 329.540 322.040 ;
        RECT 331.740 3.320 332.840 322.040 ;
        RECT 335.040 3.320 368.410 322.040 ;
        RECT 370.610 3.320 371.710 322.040 ;
        RECT 373.910 3.320 407.280 322.040 ;
        RECT 409.480 3.320 410.580 322.040 ;
        RECT 412.780 3.320 446.150 322.040 ;
        RECT 448.350 3.320 449.450 322.040 ;
        RECT 451.650 3.320 485.020 322.040 ;
        RECT 487.220 3.320 488.320 322.040 ;
        RECT 490.520 3.320 523.890 322.040 ;
        RECT 526.090 3.320 527.190 322.040 ;
        RECT 529.390 3.320 562.760 322.040 ;
        RECT 564.960 3.320 566.060 322.040 ;
        RECT 568.260 3.320 601.630 322.040 ;
        RECT 603.830 3.320 604.930 322.040 ;
        RECT 607.130 3.320 640.500 322.040 ;
        RECT 642.700 3.320 643.800 322.040 ;
        RECT 646.000 3.320 679.370 322.040 ;
        RECT 681.570 3.320 682.670 322.040 ;
        RECT 684.870 3.320 718.240 322.040 ;
        RECT 720.440 3.320 721.540 322.040 ;
        RECT 723.740 3.320 757.110 322.040 ;
        RECT 759.310 3.320 760.410 322.040 ;
        RECT 762.610 3.320 795.980 322.040 ;
        RECT 798.180 3.320 799.280 322.040 ;
        RECT 801.480 3.320 834.850 322.040 ;
        RECT 837.050 3.320 838.150 322.040 ;
        RECT 840.350 3.320 873.720 322.040 ;
        RECT 875.920 3.320 877.020 322.040 ;
        RECT 879.220 3.320 912.590 322.040 ;
        RECT 914.790 3.320 915.890 322.040 ;
        RECT 918.090 3.320 951.460 322.040 ;
        RECT 953.660 3.320 954.760 322.040 ;
        RECT 956.960 3.320 990.330 322.040 ;
        RECT 992.530 3.320 993.630 322.040 ;
        RECT 995.830 3.320 1029.200 322.040 ;
        RECT 1031.400 3.320 1032.500 322.040 ;
        RECT 1034.700 3.320 1068.070 322.040 ;
        RECT 1070.270 3.320 1071.370 322.040 ;
        RECT 1073.570 3.320 1106.940 322.040 ;
        RECT 1109.140 3.320 1110.240 322.040 ;
        RECT 1112.440 3.320 1145.810 322.040 ;
        RECT 1148.010 3.320 1149.110 322.040 ;
        RECT 1151.310 3.320 1184.680 322.040 ;
        RECT 1186.880 3.320 1187.980 322.040 ;
        RECT 1190.180 3.320 1223.550 322.040 ;
        RECT 1225.750 3.320 1226.850 322.040 ;
        RECT 1229.050 3.320 1262.420 322.040 ;
        RECT 1264.620 3.320 1265.720 322.040 ;
        RECT 1267.920 3.320 1301.290 322.040 ;
        RECT 1303.490 3.320 1304.590 322.040 ;
        RECT 1306.790 3.320 1340.160 322.040 ;
        RECT 1342.360 3.320 1343.460 322.040 ;
        RECT 1345.660 3.320 1371.300 322.040 ;
        RECT 15.260 0.090 1371.300 3.320 ;
  END
END tt_um_simple_riscv
END LIBRARY

